module AND_gate(a,b,out);
    input a, b;
    output  out
    // AND gate functionality
    assign out = a & b;

endmodule
