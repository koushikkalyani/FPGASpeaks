module EXOR_gate(a,b,out);
    input a, b;
    output  out
    // E-XOR gate functionality
    assign out = a ^ b;

endmodule
