module OR_gate(a,b,out);
    input a, b;
    output  out
    // OR gate functionality
    assign out = a | b;

endmodule

