module NOT(a,out);
   input a;
   output out;
   // NOT operation
   assign out =!a;
endmodule
